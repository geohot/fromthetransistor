
module microplexer(
  input   reg[5:0] set
  output
);

initial begin
  
end
